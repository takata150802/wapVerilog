module m0(
clk,
in0,
in1,
out0,
out1
);

input clk;
input in0;
input in1;
output out0;
output out1;
endmodule
