module m2(
clk,out
);

input clk;
output out;
endmodule
